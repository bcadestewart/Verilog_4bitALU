
module AND_Module(
    input [3:0] A,
    input [3:0] B,
    output [3:0] AND_Out
);
    assign AND_Out = A & B;
endmodule
