
module NOT_Module(
    input [3:0] A,
    output [3:0] NOT_Out
);
    assign NOT_Out = ~A;
endmodule
